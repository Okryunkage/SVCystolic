`ifndef parameter_vh
`define parameter_vh

`define clk100MHz 100_000_000
`define clk200MHz 200_000_000
`define clk300MHz 300_000_000
`define clk400MHz 400_000_000
`define clk500MHz 500_000_000

`define bitwidth5 5
`define bitwidth6 6
`define bitwidth7 7
`define bitwidth8 8

`define baud9600    9_600
`define baud19200   19_200
`define baud38400   38_400
`define baud57600   57_600
`define baud115200  115_200
`define baud230400  230_400
`define baud460800  460_800
`define baud921600  921_600

`define baud_slow   9600
`define baud_mid    115200
`define baud_fast   921600

`endif
